package apb_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "apb_txn.sv"
  `include "apb_driver.sv"
  `include "apb_monitor.sv"
  `include "apb_scoreboard.sv"
  `include "apb_env.sv"
  `include "apb_test.sv"
endpackage
